/*
IFPB
Joao Pessoa, 02 de dezembro de 2016
Aluno: Gabriel Daltro Duarte

 Disciplina System Verilog - Programa de Execelencia em Microeletronica

 Exercicio:
4) Fazer circuito que acenda os LEDs em sequência. Exemplo com 4 LEDs:

L0 L1 L2 L3

 *
      *
          *
               *
          *
      *
 *
      *
(...)


*/